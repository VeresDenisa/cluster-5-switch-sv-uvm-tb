package test_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import item_pack::*;
  import seq_pack::*;
  import base_pack::*;
  import config_pack::*;

  import env_pack::*;

  `include "src/test/test.svh"
  `include "src/test/test_no_1.svh"
  `include "src/test/test_no_2.svh"
  `include "src/test/test_no_4.svh"
  `include "src/test/test_no_5.svh"
  `include "src/test/test_no_6.svh"
  `include "src/test/test_no_7.svh"
  `include "src/test/test_no_8.svh"
  `include "src/test/test_no_9.svh"
  `include "src/test/test_no_11.svh"
  `include "src/test/test_no_12.svh"

endpackage : test_pack