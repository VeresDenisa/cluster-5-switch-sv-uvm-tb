package reset_agent_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import item_pack::*;
  import base_pack::*;
  import config_pack::*;

  `include "src/test/environment/agent_reset/reset_driver.svh"
  `include "src/test/environment/agent_reset/reset_monitor.svh"

  `include "src/test/environment/agent_reset/reset_agent.svh"
endpackage : reset_agent_pack