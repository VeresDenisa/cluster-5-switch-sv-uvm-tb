package base_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "src/test/environment/agent_base/base_agent_config.svh"

  `include "src/test/environment/agent_base/base_driver.svh"
  `include "src/test/environment/agent_base/base_monitor.svh"
  
  `include "src/test/environment/agent_base/base_agent.svh"
endpackage : base_pack