package port_agent_pack;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import item_pack::*;
  import base_pack::*;
  import config_pack::*;

  `include "src/test/environment/agent_port/port_driver.svh"
  `include "src/test/environment/agent_port/port_monitor.svh"
  `include "src/test/environment/agent_port/port_sequencer.svh"

  `include "src/test/environment/agent_port/port_agent.svh"
endpackage : port_agent_pack